//Module by Ryan Thompson
module adder_subtractor( s, op, a);


endmodule